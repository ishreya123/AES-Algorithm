//////////////////////////////////////////////////////////////////////////////////
//
// Create Date: 13.06.2025 
// Design Name: S_box
// Module Name: S_box.sv
// Project Name: AES Encryption
// Target Devices: Zed Board
// Tool Versions: Vivado 2019.1
// Description: 
// 
// Dependencies: 
// 
// Revision: v0.01
//////////////////////////////////////////////////////////////////////////////////

module S_box (a_key,c_key);
	input [7:0] a_key;
	output reg [7:0] c_key; 
	
always_comb begin : s_boxlogic
	case (a_key)

	    8'h00: c_key=8'h63;
	    8'h01: c_key=8'h7c;
	    8'h02: c_key=8'h77;
	    8'h03: c_key=8'h7b;
	    8'h04: c_key=8'hf2;
	    8'h05: c_key=8'h6b;
	    8'h06: c_key=8'h6f;
	    8'h07: c_key=8'hc5;
	    8'h08: c_key=8'h30;
	    8'h09: c_key=8'h01;
	    8'h0a: c_key=8'h67;
	    8'h0b: c_key=8'h2b;
	    8'h0c: c_key=8'hfe;
	    8'h0d: c_key=8'hd7;
	    8'h0e: c_key=8'hab;
	    8'h0f: c_key=8'h76;
	    8'h10: c_key=8'hca;
	    8'h11: c_key=8'h82;
	    8'h12: c_key=8'hc9;
	    8'h13: c_key=8'h7d;
	    8'h14: c_key=8'hfa;
	    8'h15: c_key=8'h59;
	    8'h16: c_key=8'h47;
	    8'h17: c_key=8'hf0;
	    8'h18: c_key=8'had;
	    8'h19: c_key=8'hd4;
	    8'h1a: c_key=8'ha2;
	    8'h1b: c_key=8'haf;
	    8'h1c: c_key=8'h9c;
	    8'h1d: c_key=8'ha4;
	    8'h1e: c_key=8'h72;
	    8'h1f: c_key=8'hc0;
	    8'h20: c_key=8'hb7;
	    8'h21: c_key=8'hfd;
	    8'h22: c_key=8'h93;
	    8'h23: c_key=8'h26;
	    8'h24: c_key=8'h36;
	    8'h25: c_key=8'h3f;
	    8'h26: c_key=8'hf7;
	    8'h27: c_key=8'hcc;
	    8'h28: c_key=8'h34;
	    8'h29: c_key=8'ha5;
	    8'h2a: c_key=8'he5;
	    8'h2b: c_key=8'hf1;
	    8'h2c: c_key=8'h71;
	    8'h2d: c_key=8'hd8;
	    8'h2e: c_key=8'h31;
	    8'h2f: c_key=8'h15;
	    8'h30: c_key=8'h04;
	    8'h31: c_key=8'hc7;
	    8'h32: c_key=8'h23;
	    8'h33: c_key=8'hc3;
	    8'h34: c_key=8'h18;
	    8'h35: c_key=8'h96;
 	    8'h36: c_key=8'h05;
	    8'h37: c_key=8'h9a;
	    8'h38: c_key=8'h07;
	    8'h39: c_key=8'h12;
	    8'h3a: c_key=8'h80;
	    8'h3b: c_key=8'he2;
	    8'h3c: c_key=8'heb;
	    8'h3d: c_key=8'h27;
	    8'h3e: c_key=8'hb2;
	    8'h3f: c_key=8'h75;
	    8'h40: c_key=8'h09;
	    8'h41: c_key=8'h83;
	    8'h42: c_key=8'h2c;
	    8'h43: c_key=8'h1a;
	    8'h44: c_key=8'h1b;
	    8'h45: c_key=8'h6e;
	    8'h46: c_key=8'h5a;
	    8'h47: c_key=8'ha0;
	    8'h48: c_key=8'h52;
	    8'h49: c_key=8'h3b;
	    8'h4a: c_key=8'hd6;
	    8'h4b: c_key=8'hb3;
	    8'h4c: c_key=8'h29;
	    8'h4d: c_key=8'he3;
	    8'h4e: c_key=8'h2f;
		8'h4f: c_key=8'h84;
		8'h50: c_key=8'h53;
		8'h51: c_key=8'hd1;
		8'h52: c_key=8'h00;
		8'h53: c_key=8'hed;
		8'h54: c_key=8'h20;
		8'h55: c_key=8'hfc;
		8'h56: c_key=8'hb1;
		8'h57: c_key=8'h5b;
		8'h58: c_key=8'h6a;
		8'h59: c_key=8'hcb;
		8'h5a: c_key=8'hbe;
		8'h5b: c_key=8'h39;
		8'h5c: c_key=8'h4a;
		8'h5d: c_key=8'h4c;
		8'h5e: c_key=8'h58;
		8'h5f: c_key=8'hcf;
		8'h60: c_key=8'hd0;
		8'h61: c_key=8'hef;
		8'h62: c_key=8'haa;
		8'h63: c_key=8'hfb;
		8'h64: c_key=8'h43;
		8'h65: c_key=8'h4d;
		8'h66: c_key=8'h33;
		8'h67: c_key=8'h85;
		8'h68: c_key=8'h45;
		8'h69: c_key=8'hf9;
		8'h6a: c_key=8'h02;
		8'h6b: c_key=8'h7f;
		8'h6c: c_key=8'h50;
		8'h6d: c_key=8'h3c;
		8'h6e: c_key=8'h9f;
		8'h6f: c_key=8'ha8;
		8'h70: c_key=8'h51;
		8'h71: c_key=8'ha3;
		8'h72: c_key=8'h40;
		8'h73: c_key=8'h8f;
		8'h74: c_key=8'h92;
		8'h75: c_key=8'h9d;
		8'h76: c_key=8'h38;
		8'h77: c_key=8'hf5;
		8'h78: c_key=8'hbc;
		8'h79: c_key=8'hb6;
		8'h7a: c_key=8'hda;
		8'h7b: c_key=8'h21;
		8'h7c: c_key=8'h10;
		8'h7d: c_key=8'hff;
		8'h7e: c_key=8'hf3;
		8'h7f: c_key=8'hd2;
		8'h80: c_key=8'hcd;
		8'h81: c_key=8'h0c;
		8'h82: c_key=8'h13;
		8'h83: c_key=8'hec;
		8'h84: c_key=8'h5f;
		8'h85: c_key=8'h97;
		8'h86: c_key=8'h44;
		8'h87: c_key=8'h17;
		8'h88: c_key=8'hc4;
		8'h89: c_key=8'ha7;
		8'h8a: c_key=8'h7e;
		8'h8b: c_key=8'h3d;
		8'h8c: c_key=8'h64;
		8'h8d: c_key=8'h5d;
		8'h8e: c_key=8'h19;
		8'h8f: c_key=8'h73;
		8'h90: c_key=8'h60;
		8'h91: c_key=8'h81;
		8'h92: c_key=8'h4f;
		8'h93: c_key=8'hdc;
		8'h94: c_key=8'h22;
		8'h95: c_key=8'h2a;
		8'h96: c_key=8'h90;
		8'h97: c_key=8'h88;
		8'h98: c_key=8'h46;
		8'h99: c_key=8'hee;
		8'h9a: c_key=8'hb8;
		8'h9b: c_key=8'h14;
		8'h9c: c_key=8'hde;
		8'h9d: c_key=8'h5e;
		8'h9e: c_key=8'h0b;
		8'h9f: c_key=8'hdb;
		8'ha0: c_key=8'he0;
		8'ha1: c_key=8'h32;
		8'ha2: c_key=8'h3a;
		8'ha3: c_key=8'h0a;
		8'ha4: c_key=8'h49;
		8'ha5: c_key=8'h06;
		8'ha6: c_key=8'h24;
		8'ha7: c_key=8'h5c;
		8'ha8: c_key=8'hc2;
		8'ha9: c_key=8'hd3;
		8'haa: c_key=8'hac;
		8'hab: c_key=8'h62;
		8'hac: c_key=8'h91;
		8'had: c_key=8'h95;
		8'hae: c_key=8'he4;
		8'haf: c_key=8'h79;
		8'hb0: c_key=8'he7;
		8'hb1: c_key=8'hc8;
		8'hb2: c_key=8'h37;
		8'hb3: c_key=8'h6d;
		8'hb4: c_key=8'h8d;
		8'hb5: c_key=8'hd5;
		8'hb6: c_key=8'h4e;
		8'hb7: c_key=8'ha9;
		8'hb8: c_key=8'h6c;
		8'hb9: c_key=8'h56;
		8'hba: c_key=8'hf4;
		8'hbb: c_key=8'hea;
		8'hbc: c_key=8'h65;
		8'hbd: c_key=8'h7a;
		8'hbe: c_key=8'hae;
		8'hbf: c_key=8'h08;
		8'hc0: c_key=8'hba;
		8'hc1: c_key=8'h78;
		8'hc2: c_key=8'h25;
		8'hc3: c_key=8'h2e;
		8'hc4: c_key=8'h1c;
		8'hc5: c_key=8'ha6;
		8'hc6: c_key=8'hb4;
		8'hc7: c_key=8'hc6;
		8'hc8: c_key=8'he8;
		8'hc9: c_key=8'hdd;
		8'hca: c_key=8'h74;
		8'hcb: c_key=8'h1f;
		8'hcc: c_key=8'h4b;
		8'hcd: c_key=8'hbd;
		8'hce: c_key=8'h8b;
		8'hcf: c_key=8'h8a;
		8'hd0: c_key=8'h70;
		8'hd1: c_key=8'h3e;
		8'hd2: c_key=8'hb5;
		8'hd3: c_key=8'h66;
		8'hd4: c_key=8'h48;
		8'hd5: c_key=8'h03;
		8'hd6: c_key=8'hf6;
		8'hd7: c_key=8'h0e;
		8'hd8: c_key=8'h61;
		8'hd9: c_key=8'h35;
		8'hda: c_key=8'h57;
		8'hdb: c_key=8'hb9;
		8'hdc: c_key=8'h86;
		8'hdd: c_key=8'hc1;
		8'hde: c_key=8'h1d;
		8'hdf: c_key=8'h9e;
		8'he0: c_key=8'he1;
		8'he1: c_key=8'hf8;
		8'he2: c_key=8'h98;
		8'he3: c_key=8'h11;
		8'he4: c_key=8'h69;
		8'he5: c_key=8'hd9;
		8'he6: c_key=8'h8e;
		8'he7: c_key=8'h94;
		8'he8: c_key=8'h9b;
		8'he9: c_key=8'h1e;
		8'hea: c_key=8'h87;
		8'heb: c_key=8'he9;
		8'hec: c_key=8'hce;
		8'hed: c_key=8'h55;
		8'hee: c_key=8'h28;
		8'hef: c_key=8'hdf;
		8'hf0: c_key=8'h8c;
		8'hf1: c_key=8'ha1;
		8'hf2: c_key=8'h89;
		8'hf3: c_key=8'h0d;
		8'hf4: c_key=8'hbf;
		8'hf5: c_key=8'he6;
		8'hf6: c_key=8'h42;
		8'hf7: c_key=8'h68;
		8'hf8: c_key=8'h41;
		8'hf9: c_key=8'h99;
		8'hfa: c_key=8'h2d;
		8'hfb: c_key=8'h0f;
		8'hfc: c_key=8'hb0;
		8'hfd: c_key=8'h54;
		8'hfe: c_key=8'hbb;
		8'hff: c_key=8'h16;
		//default : /* default */;
	endcase
	
end
endmodule : S_box
