class aes_transaction extends uvm_sequence_item;
  `uvm_object_utils(aes_transaction)

  function new(string name = "aes_transaction");
        super.new(name);
    endfunction
endclass
